/*
 * Order Management Module
 * Hardware-accelerated order processing and risk management
 * 
 * Features:
 * - Order state machine with 16ns latency
 * - Pre-trade risk checks
 * - Order matching engine
 * - Position tracking
 */

module order_manager #(
    parameter ORDER_WIDTH = 64,
    parameter SYMBOL_WIDTH = 32,
    parameter PRICE_WIDTH = 32,
    parameter VOLUME_WIDTH = 32,
    parameter MAX_ORDERS = 1024,
    parameter MAX_POSITIONS = 256
) (
    input  wire                     clk,
    input  wire                     rst_n,
    
    // Order input interface
    input  wire                     order_valid,
    input  wire [ORDER_WIDTH-1:0]   order_data,
    input  wire [SYMBOL_WIDTH-1:0]  order_symbol,
    input  wire [PRICE_WIDTH-1:0]   order_price,
    input  wire [VOLUME_WIDTH-1:0]  order_volume,
    input  wire                     order_side,        // 0=buy, 1=sell
    input  wire [2:0]               order_type,        // 0=market, 1=limit, 2=cancel
    input  wire [31:0]              order_id,           // Order ID input
    output wire                     order_ready,
    
    // Market data interface
    input  wire                     tick_valid,
    input  wire [SYMBOL_WIDTH-1:0]  tick_symbol,
    input  wire [PRICE_WIDTH-1:0]   tick_price,
    input  wire [PRICE_WIDTH-1:0]   tick_bid,
    input  wire [PRICE_WIDTH-1:0]   tick_ask,
    
    // Order execution output
    output reg                      exec_valid,
    output reg  [ORDER_WIDTH-1:0]   exec_order_id,
    output reg  [SYMBOL_WIDTH-1:0]  exec_symbol,
    output reg  [PRICE_WIDTH-1:0]   exec_price,
    output reg  [VOLUME_WIDTH-1:0]  exec_volume,
    output reg                      exec_side,
    output reg  [63:0]              exec_timestamp,
    
    // Position updates
    output reg                      pos_update_valid,
    output reg  [SYMBOL_WIDTH-1:0]  pos_symbol,
    output reg  [VOLUME_WIDTH-1:0]  pos_quantity,
    output reg                      pos_side,
    
    // Risk management interface
    input  wire [PRICE_WIDTH-1:0]   risk_position_limit,
    input  wire [PRICE_WIDTH-1:0]   risk_max_order_size,
    input  wire                     risk_enabled,
    output wire                     risk_violation,
    
    // Statistics
    output wire [31:0]              orders_processed,
    output wire [31:0]              orders_filled,
    output wire [31:0]              orders_rejected,
    output wire [15:0]              active_orders,
    
    // Additional outputs
    output wire [31:0]              risk_code,          // Risk code output
    output wire [31:0]              execution_status,   // Execution status output
    output wire [31:0]              position_pnl       // Position PnL output
);

// Internal registers
reg [31:0] order_counter;
reg [31:0] fill_counter;
reg [31:0] reject_counter;
reg [15:0] active_order_count;

// Loop variable for initialization
integer i;

// Order state machine
localparam ORDER_IDLE = 3'b000;
localparam ORDER_VALIDATE = 3'b001;
localparam ORDER_RISK_CHECK = 3'b010;
localparam ORDER_MATCH = 3'b011;
localparam ORDER_EXECUTE = 3'b100;
localparam ORDER_REJECT = 3'b101;
localparam ORDER_COMPLETE = 3'b110;

reg [2:0] order_state;
reg [2:0] next_order_state;

// Order storage (simplified - in real implementation would use CAM/TCAM)
reg [ORDER_WIDTH-1:0]   order_memory [0:MAX_ORDERS-1];
reg [SYMBOL_WIDTH-1:0]  order_symbols [0:MAX_ORDERS-1];
reg [PRICE_WIDTH-1:0]   order_prices [0:MAX_ORDERS-1];
reg [VOLUME_WIDTH-1:0]  order_volumes [0:MAX_ORDERS-1];
reg                     order_sides [0:MAX_ORDERS-1];
reg [2:0]               order_types [0:MAX_ORDERS-1];
reg                     order_valid_flags [0:MAX_ORDERS-1];
reg [9:0]               order_write_ptr;
reg [9:0]               order_read_ptr;

// Position tracking
reg [VOLUME_WIDTH-1:0]  positions [0:MAX_POSITIONS-1];
reg [SYMBOL_WIDTH-1:0]  position_symbols [0:MAX_POSITIONS-1];
reg [7:0]               position_count;

// Current order being processed
reg [ORDER_WIDTH-1:0]   current_order;
reg [SYMBOL_WIDTH-1:0]  current_symbol;
reg [PRICE_WIDTH-1:0]   current_price;
reg [VOLUME_WIDTH-1:0]  current_volume;
reg                     current_side;
reg [2:0]               current_type;

// Risk check results
wire risk_position_ok;
wire risk_size_ok;
wire risk_all_ok;

// Matching engine
wire match_found;
wire [PRICE_WIDTH-1:0] match_price;
wire [VOLUME_WIDTH-1:0] match_volume;

// Pipeline timing
reg [3:0] pipeline_counter;

// Statistics outputs
assign orders_processed = order_counter;
assign orders_filled = fill_counter;
assign orders_rejected = reject_counter;
assign active_orders = active_order_count;

// Order ready signal
assign order_ready = (order_state == ORDER_IDLE) || (order_state == ORDER_COMPLETE);

// Risk violation output
assign risk_violation = risk_violation_sticky;

// Risk code logic
assign risk_code = !risk_position_ok ? 32'd1 :
                   !risk_size_ok     ? 32'd2 : 32'd0;

// Execution status logic
assign execution_status = (order_state == ORDER_EXECUTE) ? 32'd1 :
                         (order_state == ORDER_REJECT)  ? 32'd2 : 32'd0;

// Position PnL logic (placeholder)
assign position_pnl = 32'd0;

// Sticky signals for testbench visibility
reg exec_valid_sticky;
reg pos_update_valid_sticky;
reg risk_violation_sticky;

// Main state machine
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        order_state <= ORDER_IDLE;
        order_counter <= 32'b0;
        fill_counter <= 32'b0;
        reject_counter <= 32'b0;
        active_order_count <= 16'b0;
        order_write_ptr <= 10'b0;
        order_read_ptr <= 10'b0;
        position_count <= 8'b0;
        pipeline_counter <= 4'b0;
        
        exec_valid <= 1'b0;
        pos_update_valid <= 1'b0;
        exec_valid_sticky <= 1'b0;
        pos_update_valid_sticky <= 1'b0;
        risk_violation_sticky <= 1'b0;
        
        // Initialize order memory
        for (i = 0; i < MAX_ORDERS; i = i + 1) begin
            order_valid_flags[i] <= 1'b0;
        end
        
    end else begin
        case (order_state)
            ORDER_IDLE: begin
                exec_valid <= 1'b0;
                pos_update_valid <= 1'b0;
                pipeline_counter <= 4'b0;
                
                if (order_valid) begin
                    // Capture new order
                    current_order <= {32'b0, order_id};
                    current_symbol <= order_symbol;
                    current_price <= order_price;
                    current_volume <= order_volume;
                    current_side <= order_side;
                    current_type <= order_type;
                    
                    order_state <= ORDER_VALIDATE;
                    pipeline_counter <= 4'b1;
                end
            end
            
            ORDER_VALIDATE: begin
                pipeline_counter <= pipeline_counter + 1;
                
                // Basic validation (1 clock cycle)
                if (current_volume == 0 || current_price == 0) begin
                    order_state <= ORDER_REJECT;
                end else begin
                    order_state <= ORDER_RISK_CHECK;
                end
            end
            
            ORDER_RISK_CHECK: begin
                pipeline_counter <= pipeline_counter + 1;
                
                // Risk checks (1 clock cycle)
                if (risk_enabled && !risk_all_ok) begin
                    order_state <= ORDER_REJECT;
                end else begin
                    order_state <= ORDER_MATCH;
                end
            end
            
            ORDER_MATCH: begin
                pipeline_counter <= pipeline_counter + 1;
                
                // Order matching logic (1 clock cycle)
                if (current_type == 3'b000) begin  // Market order
                    order_state <= ORDER_EXECUTE;
                end else if (current_type == 3'b001) begin  // Limit order
                    if (match_found) begin
                        order_state <= ORDER_EXECUTE;
                    end else begin
                        // Store order for later matching
                        order_memory[order_write_ptr] <= current_order;
                        order_symbols[order_write_ptr] <= current_symbol;
                        order_prices[order_write_ptr] <= current_price;
                        order_volumes[order_write_ptr] <= current_volume;
                        order_sides[order_write_ptr] <= current_side;
                        order_types[order_write_ptr] <= current_type;
                        order_valid_flags[order_write_ptr] <= 1'b1;
                        
                        order_write_ptr <= order_write_ptr + 1;
                        active_order_count <= active_order_count + 1;
                        
                        order_state <= ORDER_COMPLETE;
                    end
                end else begin  // Cancel order
                    // Cancel logic would go here
                    order_state <= ORDER_COMPLETE;
                end
            end
            
            ORDER_EXECUTE: begin
                pipeline_counter <= pipeline_counter + 1;
                
                // Execute order (1 clock cycle)
                exec_valid <= 1'b1;
                exec_order_id <= current_order;
                exec_symbol <= current_symbol;
                exec_price <= (current_type == 3'b000) ? 
                             (current_side ? tick_ask : tick_bid) : current_price;
                exec_volume <= current_volume;
                exec_side <= current_side;
                exec_timestamp <= $time;
                
                // Update position
                pos_update_valid <= 1'b1;
                pos_symbol <= current_symbol;
                pos_quantity <= current_volume;
                pos_side <= current_side;
                
                fill_counter <= fill_counter + 1;
                order_state <= ORDER_COMPLETE;
            end
            
            ORDER_REJECT: begin
                reject_counter <= reject_counter + 1;
                order_state <= ORDER_COMPLETE;
            end
            
            ORDER_COMPLETE: begin
                order_counter <= order_counter + 1;
                order_state <= ORDER_IDLE;
            end
            
            default: begin
                order_state <= ORDER_IDLE;
            end
        endcase
    end
end

// Risk management logic
assign risk_position_ok = !risk_enabled || (current_volume <= risk_position_limit);
assign risk_size_ok = !risk_enabled || (current_volume <= risk_max_order_size);
assign risk_all_ok = risk_position_ok && risk_size_ok;

// Simple matching engine (combinational logic)
assign match_found = (current_type == 3'b001) && tick_valid && 
                    (current_symbol == tick_symbol) &&
                    ((current_side == 1'b0 && current_price >= tick_ask) ||
                     (current_side == 1'b1 && current_price <= tick_bid));

assign match_price = current_side ? tick_bid : tick_ask;
assign match_volume = current_volume;  // Simplified - assume full fill

// Position management
integer pos_idx;
reg position_found;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        // Initialize positions
        integer j;
        for (j = 0; j < MAX_POSITIONS; j = j + 1) begin
            positions[j] <= {VOLUME_WIDTH{1'b0}};
            position_symbols[j] <= {SYMBOL_WIDTH{1'b0}};
        end
    end else if (pos_update_valid) begin
        // Update position
        position_found = 1'b0;
        
        for (pos_idx = 0; pos_idx < position_count; pos_idx = pos_idx + 1) begin
            if (position_symbols[pos_idx] == pos_symbol) begin
                if (pos_side == 1'b0) begin  // Buy
                    positions[pos_idx] <= positions[pos_idx] + pos_quantity;
                end else begin  // Sell
                    positions[pos_idx] <= positions[pos_idx] - pos_quantity;
                end
                position_found = 1'b1;
            end
        end
        
        // Add new position if symbol not found
        if (!position_found && position_count < MAX_POSITIONS) begin
            position_symbols[position_count] <= pos_symbol;
            positions[position_count] <= pos_side ? -pos_quantity : pos_quantity;
            position_count <= position_count + 1;
        end
    end
end

endmodule
